`define WT_DCACHE
